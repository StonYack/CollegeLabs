// Lab3Nios.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module Lab3Nios (
		input  wire        clk_clk,         //      clk.clk
		output wire [20:0] hex_export,      //      hex.export
		input  wire [9:0]  switches_export  // switches.export
	);

	wire         lab3nios_debug_reset_request_reset;                          // Lab3Nios:debug_reset_request -> rst_controller:reset_in0
	wire  [31:0] lab3nios_data_master_readdata;                               // mm_interconnect_0:Lab3Nios_data_master_readdata -> Lab3Nios:d_readdata
	wire         lab3nios_data_master_waitrequest;                            // mm_interconnect_0:Lab3Nios_data_master_waitrequest -> Lab3Nios:d_waitrequest
	wire         lab3nios_data_master_debugaccess;                            // Lab3Nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Lab3Nios_data_master_debugaccess
	wire  [13:0] lab3nios_data_master_address;                                // Lab3Nios:d_address -> mm_interconnect_0:Lab3Nios_data_master_address
	wire   [3:0] lab3nios_data_master_byteenable;                             // Lab3Nios:d_byteenable -> mm_interconnect_0:Lab3Nios_data_master_byteenable
	wire         lab3nios_data_master_read;                                   // Lab3Nios:d_read -> mm_interconnect_0:Lab3Nios_data_master_read
	wire         lab3nios_data_master_readdatavalid;                          // mm_interconnect_0:Lab3Nios_data_master_readdatavalid -> Lab3Nios:d_readdatavalid
	wire         lab3nios_data_master_write;                                  // Lab3Nios:d_write -> mm_interconnect_0:Lab3Nios_data_master_write
	wire  [31:0] lab3nios_data_master_writedata;                              // Lab3Nios:d_writedata -> mm_interconnect_0:Lab3Nios_data_master_writedata
	wire  [31:0] lab3nios_instruction_master_readdata;                        // mm_interconnect_0:Lab3Nios_instruction_master_readdata -> Lab3Nios:i_readdata
	wire         lab3nios_instruction_master_waitrequest;                     // mm_interconnect_0:Lab3Nios_instruction_master_waitrequest -> Lab3Nios:i_waitrequest
	wire  [13:0] lab3nios_instruction_master_address;                         // Lab3Nios:i_address -> mm_interconnect_0:Lab3Nios_instruction_master_address
	wire         lab3nios_instruction_master_read;                            // Lab3Nios:i_read -> mm_interconnect_0:Lab3Nios_instruction_master_read
	wire         lab3nios_instruction_master_readdatavalid;                   // mm_interconnect_0:Lab3Nios_instruction_master_readdatavalid -> Lab3Nios:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_lab3nios_debug_mem_slave_readdata;         // Lab3Nios:debug_mem_slave_readdata -> mm_interconnect_0:Lab3Nios_debug_mem_slave_readdata
	wire         mm_interconnect_0_lab3nios_debug_mem_slave_waitrequest;      // Lab3Nios:debug_mem_slave_waitrequest -> mm_interconnect_0:Lab3Nios_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_lab3nios_debug_mem_slave_debugaccess;      // mm_interconnect_0:Lab3Nios_debug_mem_slave_debugaccess -> Lab3Nios:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_lab3nios_debug_mem_slave_address;          // mm_interconnect_0:Lab3Nios_debug_mem_slave_address -> Lab3Nios:debug_mem_slave_address
	wire         mm_interconnect_0_lab3nios_debug_mem_slave_read;             // mm_interconnect_0:Lab3Nios_debug_mem_slave_read -> Lab3Nios:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_lab3nios_debug_mem_slave_byteenable;       // mm_interconnect_0:Lab3Nios_debug_mem_slave_byteenable -> Lab3Nios:debug_mem_slave_byteenable
	wire         mm_interconnect_0_lab3nios_debug_mem_slave_write;            // mm_interconnect_0:Lab3Nios_debug_mem_slave_write -> Lab3Nios:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_lab3nios_debug_mem_slave_writedata;        // mm_interconnect_0:Lab3Nios_debug_mem_slave_writedata -> Lab3Nios:debug_mem_slave_writedata
	wire         mm_interconnect_0_memory_s1_chipselect;                      // mm_interconnect_0:Memory_s1_chipselect -> Memory:chipselect
	wire  [31:0] mm_interconnect_0_memory_s1_readdata;                        // Memory:readdata -> mm_interconnect_0:Memory_s1_readdata
	wire   [9:0] mm_interconnect_0_memory_s1_address;                         // mm_interconnect_0:Memory_s1_address -> Memory:address
	wire   [3:0] mm_interconnect_0_memory_s1_byteenable;                      // mm_interconnect_0:Memory_s1_byteenable -> Memory:byteenable
	wire         mm_interconnect_0_memory_s1_write;                           // mm_interconnect_0:Memory_s1_write -> Memory:write
	wire  [31:0] mm_interconnect_0_memory_s1_writedata;                       // mm_interconnect_0:Memory_s1_writedata -> Memory:writedata
	wire         mm_interconnect_0_memory_s1_clken;                           // mm_interconnect_0:Memory_s1_clken -> Memory:clken
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                      // Switches:readdata -> mm_interconnect_0:Switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                       // mm_interconnect_0:Switches_s1_address -> Switches:address
	wire         mm_interconnect_0_hex_s1_chipselect;                         // mm_interconnect_0:Hex_s1_chipselect -> Hex:chipselect
	wire  [31:0] mm_interconnect_0_hex_s1_readdata;                           // Hex:readdata -> mm_interconnect_0:Hex_s1_readdata
	wire   [1:0] mm_interconnect_0_hex_s1_address;                            // mm_interconnect_0:Hex_s1_address -> Hex:address
	wire         mm_interconnect_0_hex_s1_write;                              // mm_interconnect_0:Hex_s1_write -> Hex:write_n
	wire  [31:0] mm_interconnect_0_hex_s1_writedata;                          // mm_interconnect_0:Hex_s1_writedata -> Hex:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] lab3nios_irq_irq;                                            // irq_mapper:sender_irq -> Lab3Nios:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [Hex:reset_n, Lab3Nios:reset_n, Memory:reset, Switches:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:Lab3Nios_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [Lab3Nios:reset_req, Memory:reset_req, rst_translator:reset_req_in]

	Lab3Nios_Hex hex (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_hex_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex_s1_readdata),   //                    .readdata
		.out_port   (hex_export)                           // external_connection.export
	);

	Lab3Nios_Lab3Nios lab3nios (
		.clk                                 (clk_clk),                                                //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (lab3nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (lab3nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (lab3nios_data_master_read),                              //                          .read
		.d_readdata                          (lab3nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (lab3nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (lab3nios_data_master_write),                             //                          .write
		.d_writedata                         (lab3nios_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (lab3nios_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (lab3nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (lab3nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (lab3nios_instruction_master_read),                       //                          .read
		.i_readdata                          (lab3nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (lab3nios_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (lab3nios_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (lab3nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (lab3nios_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_lab3nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_lab3nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_lab3nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_lab3nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_lab3nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_lab3nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_lab3nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_lab3nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                        // custom_instruction_master.readra
	);

	Lab3Nios_Memory memory (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	Lab3Nios_Switches switches (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	Lab3Nios_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	Lab3Nios_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                              (clk_clk),                                                     //                            clk_0_clk.clk
		.Lab3Nios_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // Lab3Nios_reset_reset_bridge_in_reset.reset
		.Lab3Nios_data_master_address               (lab3nios_data_master_address),                                //                 Lab3Nios_data_master.address
		.Lab3Nios_data_master_waitrequest           (lab3nios_data_master_waitrequest),                            //                                     .waitrequest
		.Lab3Nios_data_master_byteenable            (lab3nios_data_master_byteenable),                             //                                     .byteenable
		.Lab3Nios_data_master_read                  (lab3nios_data_master_read),                                   //                                     .read
		.Lab3Nios_data_master_readdata              (lab3nios_data_master_readdata),                               //                                     .readdata
		.Lab3Nios_data_master_readdatavalid         (lab3nios_data_master_readdatavalid),                          //                                     .readdatavalid
		.Lab3Nios_data_master_write                 (lab3nios_data_master_write),                                  //                                     .write
		.Lab3Nios_data_master_writedata             (lab3nios_data_master_writedata),                              //                                     .writedata
		.Lab3Nios_data_master_debugaccess           (lab3nios_data_master_debugaccess),                            //                                     .debugaccess
		.Lab3Nios_instruction_master_address        (lab3nios_instruction_master_address),                         //          Lab3Nios_instruction_master.address
		.Lab3Nios_instruction_master_waitrequest    (lab3nios_instruction_master_waitrequest),                     //                                     .waitrequest
		.Lab3Nios_instruction_master_read           (lab3nios_instruction_master_read),                            //                                     .read
		.Lab3Nios_instruction_master_readdata       (lab3nios_instruction_master_readdata),                        //                                     .readdata
		.Lab3Nios_instruction_master_readdatavalid  (lab3nios_instruction_master_readdatavalid),                   //                                     .readdatavalid
		.Hex_s1_address                             (mm_interconnect_0_hex_s1_address),                            //                               Hex_s1.address
		.Hex_s1_write                               (mm_interconnect_0_hex_s1_write),                              //                                     .write
		.Hex_s1_readdata                            (mm_interconnect_0_hex_s1_readdata),                           //                                     .readdata
		.Hex_s1_writedata                           (mm_interconnect_0_hex_s1_writedata),                          //                                     .writedata
		.Hex_s1_chipselect                          (mm_interconnect_0_hex_s1_chipselect),                         //                                     .chipselect
		.jtag_uart_0_avalon_jtag_slave_address      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //        jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                     .write
		.jtag_uart_0_avalon_jtag_slave_read         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                     .read
		.jtag_uart_0_avalon_jtag_slave_readdata     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                     .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                     .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                     .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                     .chipselect
		.Lab3Nios_debug_mem_slave_address           (mm_interconnect_0_lab3nios_debug_mem_slave_address),          //             Lab3Nios_debug_mem_slave.address
		.Lab3Nios_debug_mem_slave_write             (mm_interconnect_0_lab3nios_debug_mem_slave_write),            //                                     .write
		.Lab3Nios_debug_mem_slave_read              (mm_interconnect_0_lab3nios_debug_mem_slave_read),             //                                     .read
		.Lab3Nios_debug_mem_slave_readdata          (mm_interconnect_0_lab3nios_debug_mem_slave_readdata),         //                                     .readdata
		.Lab3Nios_debug_mem_slave_writedata         (mm_interconnect_0_lab3nios_debug_mem_slave_writedata),        //                                     .writedata
		.Lab3Nios_debug_mem_slave_byteenable        (mm_interconnect_0_lab3nios_debug_mem_slave_byteenable),       //                                     .byteenable
		.Lab3Nios_debug_mem_slave_waitrequest       (mm_interconnect_0_lab3nios_debug_mem_slave_waitrequest),      //                                     .waitrequest
		.Lab3Nios_debug_mem_slave_debugaccess       (mm_interconnect_0_lab3nios_debug_mem_slave_debugaccess),      //                                     .debugaccess
		.Memory_s1_address                          (mm_interconnect_0_memory_s1_address),                         //                            Memory_s1.address
		.Memory_s1_write                            (mm_interconnect_0_memory_s1_write),                           //                                     .write
		.Memory_s1_readdata                         (mm_interconnect_0_memory_s1_readdata),                        //                                     .readdata
		.Memory_s1_writedata                        (mm_interconnect_0_memory_s1_writedata),                       //                                     .writedata
		.Memory_s1_byteenable                       (mm_interconnect_0_memory_s1_byteenable),                      //                                     .byteenable
		.Memory_s1_chipselect                       (mm_interconnect_0_memory_s1_chipselect),                      //                                     .chipselect
		.Memory_s1_clken                            (mm_interconnect_0_memory_s1_clken),                           //                                     .clken
		.Switches_s1_address                        (mm_interconnect_0_switches_s1_address),                       //                          Switches_s1.address
		.Switches_s1_readdata                       (mm_interconnect_0_switches_s1_readdata)                       //                                     .readdata
	);

	Lab3Nios_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (lab3nios_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (lab3nios_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
