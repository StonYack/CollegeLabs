// FreeRTOS.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module FreeRTOS (
		input  wire        clk_clk,          //        clk.clk
		output wire [6:0]  hex_0_export,     //      hex_0.export
		output wire [5:0]  piezo_0_export,   //    piezo_0.export
		output wire        sdram_clk_clk,    //  sdram_clk.clk
		output wire [12:0] sdram_wire_addr,  // sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,    //           .ba
		output wire        sdram_wire_cas_n, //           .cas_n
		output wire        sdram_wire_cke,   //           .cke
		output wire        sdram_wire_cs_n,  //           .cs_n
		inout  wire [15:0] sdram_wire_dq,    //           .dq
		output wire [1:0]  sdram_wire_dqm,   //           .dqm
		output wire        sdram_wire_ras_n, //           .ras_n
		output wire        sdram_wire_we_n,  //           .we_n
		output wire [5:0]  servo_0_export,   //    servo_0.export
		output wire [5:0]  servo_1_export,   //    servo_1.export
		input  wire [3:0]  sw_0_export       //       sw_0.export
	);

	wire         clock_sys_clk_clk;                                           // clock:sys_clk_clk -> [FreeRTOSNios:clk, Hex_0:clk, Piezo_0:clk, SW_0:clk, Servo_0:clk, Servo_1:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:clock_sys_clk_clk, rst_controller:clk, sdram:clk, sys_clk:clk, timer_0:clk, timer_1:clk, timer_2:clk]
	wire         freertosnios_debug_reset_request_reset;                      // FreeRTOSNios:debug_reset_request -> [clock:ref_reset_reset, rst_controller:reset_in0]
	wire  [31:0] freertosnios_data_master_readdata;                           // mm_interconnect_0:FreeRTOSNios_data_master_readdata -> FreeRTOSNios:d_readdata
	wire         freertosnios_data_master_waitrequest;                        // mm_interconnect_0:FreeRTOSNios_data_master_waitrequest -> FreeRTOSNios:d_waitrequest
	wire         freertosnios_data_master_debugaccess;                        // FreeRTOSNios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:FreeRTOSNios_data_master_debugaccess
	wire  [27:0] freertosnios_data_master_address;                            // FreeRTOSNios:d_address -> mm_interconnect_0:FreeRTOSNios_data_master_address
	wire   [3:0] freertosnios_data_master_byteenable;                         // FreeRTOSNios:d_byteenable -> mm_interconnect_0:FreeRTOSNios_data_master_byteenable
	wire         freertosnios_data_master_read;                               // FreeRTOSNios:d_read -> mm_interconnect_0:FreeRTOSNios_data_master_read
	wire         freertosnios_data_master_readdatavalid;                      // mm_interconnect_0:FreeRTOSNios_data_master_readdatavalid -> FreeRTOSNios:d_readdatavalid
	wire         freertosnios_data_master_write;                              // FreeRTOSNios:d_write -> mm_interconnect_0:FreeRTOSNios_data_master_write
	wire  [31:0] freertosnios_data_master_writedata;                          // FreeRTOSNios:d_writedata -> mm_interconnect_0:FreeRTOSNios_data_master_writedata
	wire  [31:0] freertosnios_instruction_master_readdata;                    // mm_interconnect_0:FreeRTOSNios_instruction_master_readdata -> FreeRTOSNios:i_readdata
	wire         freertosnios_instruction_master_waitrequest;                 // mm_interconnect_0:FreeRTOSNios_instruction_master_waitrequest -> FreeRTOSNios:i_waitrequest
	wire  [27:0] freertosnios_instruction_master_address;                     // FreeRTOSNios:i_address -> mm_interconnect_0:FreeRTOSNios_instruction_master_address
	wire         freertosnios_instruction_master_read;                        // FreeRTOSNios:i_read -> mm_interconnect_0:FreeRTOSNios_instruction_master_read
	wire         freertosnios_instruction_master_readdatavalid;               // mm_interconnect_0:FreeRTOSNios_instruction_master_readdatavalid -> FreeRTOSNios:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_hex_0_avalon_slave_0_chipselect;           // mm_interconnect_0:Hex_0_avalon_slave_0_chipselect -> Hex_0:chipselect
	wire  [31:0] mm_interconnect_0_hex_0_avalon_slave_0_readdata;             // Hex_0:readdata -> mm_interconnect_0:Hex_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_hex_0_avalon_slave_0_address;              // mm_interconnect_0:Hex_0_avalon_slave_0_address -> Hex_0:address
	wire         mm_interconnect_0_hex_0_avalon_slave_0_write;                // mm_interconnect_0:Hex_0_avalon_slave_0_write -> Hex_0:write_n
	wire  [31:0] mm_interconnect_0_hex_0_avalon_slave_0_writedata;            // mm_interconnect_0:Hex_0_avalon_slave_0_writedata -> Hex_0:writedata
	wire  [31:0] mm_interconnect_0_sw_0_avalon_slave_0_readdata;              // SW_0:readdata -> mm_interconnect_0:SW_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_sw_0_avalon_slave_0_address;               // mm_interconnect_0:SW_0_avalon_slave_0_address -> SW_0:address
	wire         mm_interconnect_0_piezo_0_avalon_slave_0_chipselect;         // mm_interconnect_0:Piezo_0_avalon_slave_0_chipselect -> Piezo_0:chipselect
	wire  [31:0] mm_interconnect_0_piezo_0_avalon_slave_0_readdata;           // Piezo_0:readdata -> mm_interconnect_0:Piezo_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_piezo_0_avalon_slave_0_address;            // mm_interconnect_0:Piezo_0_avalon_slave_0_address -> Piezo_0:address
	wire         mm_interconnect_0_piezo_0_avalon_slave_0_write;              // mm_interconnect_0:Piezo_0_avalon_slave_0_write -> Piezo_0:write_n
	wire  [31:0] mm_interconnect_0_piezo_0_avalon_slave_0_writedata;          // mm_interconnect_0:Piezo_0_avalon_slave_0_writedata -> Piezo_0:writedata
	wire         mm_interconnect_0_servo_0_avalon_slave_0_chipselect;         // mm_interconnect_0:Servo_0_avalon_slave_0_chipselect -> Servo_0:chipselect
	wire  [31:0] mm_interconnect_0_servo_0_avalon_slave_0_readdata;           // Servo_0:readdata -> mm_interconnect_0:Servo_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_servo_0_avalon_slave_0_address;            // mm_interconnect_0:Servo_0_avalon_slave_0_address -> Servo_0:address
	wire         mm_interconnect_0_servo_0_avalon_slave_0_write;              // mm_interconnect_0:Servo_0_avalon_slave_0_write -> Servo_0:write_n
	wire  [31:0] mm_interconnect_0_servo_0_avalon_slave_0_writedata;          // mm_interconnect_0:Servo_0_avalon_slave_0_writedata -> Servo_0:writedata
	wire         mm_interconnect_0_servo_1_avalon_slave_0_chipselect;         // mm_interconnect_0:Servo_1_avalon_slave_0_chipselect -> Servo_1:chipselect
	wire  [31:0] mm_interconnect_0_servo_1_avalon_slave_0_readdata;           // Servo_1:readdata -> mm_interconnect_0:Servo_1_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_servo_1_avalon_slave_0_address;            // mm_interconnect_0:Servo_1_avalon_slave_0_address -> Servo_1:address
	wire         mm_interconnect_0_servo_1_avalon_slave_0_write;              // mm_interconnect_0:Servo_1_avalon_slave_0_write -> Servo_1:write_n
	wire  [31:0] mm_interconnect_0_servo_1_avalon_slave_0_writedata;          // mm_interconnect_0:Servo_1_avalon_slave_0_writedata -> Servo_1:writedata
	wire  [31:0] mm_interconnect_0_freertosnios_debug_mem_slave_readdata;     // FreeRTOSNios:debug_mem_slave_readdata -> mm_interconnect_0:FreeRTOSNios_debug_mem_slave_readdata
	wire         mm_interconnect_0_freertosnios_debug_mem_slave_waitrequest;  // FreeRTOSNios:debug_mem_slave_waitrequest -> mm_interconnect_0:FreeRTOSNios_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_freertosnios_debug_mem_slave_debugaccess;  // mm_interconnect_0:FreeRTOSNios_debug_mem_slave_debugaccess -> FreeRTOSNios:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_freertosnios_debug_mem_slave_address;      // mm_interconnect_0:FreeRTOSNios_debug_mem_slave_address -> FreeRTOSNios:debug_mem_slave_address
	wire         mm_interconnect_0_freertosnios_debug_mem_slave_read;         // mm_interconnect_0:FreeRTOSNios_debug_mem_slave_read -> FreeRTOSNios:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_freertosnios_debug_mem_slave_byteenable;   // mm_interconnect_0:FreeRTOSNios_debug_mem_slave_byteenable -> FreeRTOSNios:debug_mem_slave_byteenable
	wire         mm_interconnect_0_freertosnios_debug_mem_slave_write;        // mm_interconnect_0:FreeRTOSNios_debug_mem_slave_write -> FreeRTOSNios:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_freertosnios_debug_mem_slave_writedata;    // mm_interconnect_0:FreeRTOSNios_debug_mem_slave_writedata -> FreeRTOSNios:debug_mem_slave_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_sys_clk_s1_chipselect;                     // mm_interconnect_0:sys_clk_s1_chipselect -> sys_clk:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_s1_readdata;                       // sys_clk:readdata -> mm_interconnect_0:sys_clk_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_s1_address;                        // mm_interconnect_0:sys_clk_s1_address -> sys_clk:address
	wire         mm_interconnect_0_sys_clk_s1_write;                          // mm_interconnect_0:sys_clk_s1_write -> sys_clk:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_s1_writedata;                      // mm_interconnect_0:sys_clk_s1_writedata -> sys_clk:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                     // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                       // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                        // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                          // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                      // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         mm_interconnect_0_timer_2_s1_chipselect;                     // mm_interconnect_0:timer_2_s1_chipselect -> timer_2:chipselect
	wire  [15:0] mm_interconnect_0_timer_2_s1_readdata;                       // timer_2:readdata -> mm_interconnect_0:timer_2_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_2_s1_address;                        // mm_interconnect_0:timer_2_s1_address -> timer_2:address
	wire         mm_interconnect_0_timer_2_s1_write;                          // mm_interconnect_0:timer_2_s1_write -> timer_2:write_n
	wire  [15:0] mm_interconnect_0_timer_2_s1_writedata;                      // mm_interconnect_0:timer_2_s1_writedata -> timer_2:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // sys_clk:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // timer_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // timer_1:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                    // timer_2:irq -> irq_mapper:receiver4_irq
	wire  [31:0] freertosnios_irq_irq;                                        // irq_mapper:sender_irq -> FreeRTOSNios:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [FreeRTOSNios:reset_n, Hex_0:reset_n, Piezo_0:reset_n, SW_0:reset_n, Servo_0:reset_n, Servo_1:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:FreeRTOSNios_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, sys_clk:reset_n, timer_0:reset_n, timer_1:reset_n, timer_2:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [FreeRTOSNios:reset_req, rst_translator:reset_req_in]

	FreeRTOS_FreeRTOSNios freertosnios (
		.clk                                 (clock_sys_clk_clk),                                          //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (freertosnios_data_master_address),                           //               data_master.address
		.d_byteenable                        (freertosnios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (freertosnios_data_master_read),                              //                          .read
		.d_readdata                          (freertosnios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (freertosnios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (freertosnios_data_master_write),                             //                          .write
		.d_writedata                         (freertosnios_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (freertosnios_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (freertosnios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (freertosnios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (freertosnios_instruction_master_read),                       //                          .read
		.i_readdata                          (freertosnios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (freertosnios_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (freertosnios_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (freertosnios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (freertosnios_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_freertosnios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_freertosnios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_freertosnios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_freertosnios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_freertosnios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_freertosnios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_freertosnios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_freertosnios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	Hex hex_0 (
		.address    (mm_interconnect_0_hex_0_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_hex_0_avalon_slave_0_chipselect), //               .chipselect
		.write_n    (~mm_interconnect_0_hex_0_avalon_slave_0_write),     //               .write_n
		.writedata  (mm_interconnect_0_hex_0_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_hex_0_avalon_slave_0_readdata),   //               .readdata
		.clk        (clock_sys_clk_clk),                                 //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //          reset.reset_n
		.out_port   (hex_0_export)                                       //    conduit_end.export
	);

	Piezo piezo_0 (
		.address    (mm_interconnect_0_piezo_0_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_piezo_0_avalon_slave_0_chipselect), //               .chipselect
		.write_n    (~mm_interconnect_0_piezo_0_avalon_slave_0_write),     //               .write_n
		.writedata  (mm_interconnect_0_piezo_0_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_piezo_0_avalon_slave_0_readdata),   //               .readdata
		.clk        (clock_sys_clk_clk),                                   //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //          reset.reset_n
		.out_port   (piezo_0_export)                                       //    conduit_end.export
	);

	SW sw_0 (
		.address  (mm_interconnect_0_sw_0_avalon_slave_0_address),  // avalon_slave_0.address
		.readdata (mm_interconnect_0_sw_0_avalon_slave_0_readdata), //               .readdata
		.clk      (clock_sys_clk_clk),                              //          clock.clk
		.reset_n  (~rst_controller_reset_out_reset),                //          reset.reset_n
		.SW_in    (sw_0_export)                                     //    conduit_end.export
	);

	Servo servo_0 (
		.address    (mm_interconnect_0_servo_0_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_servo_0_avalon_slave_0_chipselect), //               .chipselect
		.write_n    (~mm_interconnect_0_servo_0_avalon_slave_0_write),     //               .write_n
		.writedata  (mm_interconnect_0_servo_0_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_servo_0_avalon_slave_0_readdata),   //               .readdata
		.clk        (clock_sys_clk_clk),                                   //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //          reset.reset_n
		.out_port   (servo_0_export)                                       //    conduit_end.export
	);

	Servo servo_1 (
		.address    (mm_interconnect_0_servo_1_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_servo_1_avalon_slave_0_chipselect), //               .chipselect
		.write_n    (~mm_interconnect_0_servo_1_avalon_slave_0_write),     //               .write_n
		.writedata  (mm_interconnect_0_servo_1_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_servo_1_avalon_slave_0_readdata),   //               .readdata
		.clk        (clock_sys_clk_clk),                                   //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                     //          reset.reset_n
		.out_port   (servo_1_export)                                       //    conduit_end.export
	);

	FreeRTOS_clock clock (
		.ref_clk_clk        (clk_clk),                                //      ref_clk.clk
		.ref_reset_reset    (freertosnios_debug_reset_request_reset), //    ref_reset.reset
		.sys_clk_clk        (clock_sys_clk_clk),                      //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                          //    sdram_clk.clk
		.reset_source_reset ()                                        // reset_source.reset
	);

	FreeRTOS_jtag_uart_0 jtag_uart_0 (
		.clk            (clock_sys_clk_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	FreeRTOS_sdram sdram (
		.clk            (clock_sys_clk_clk),                        //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	FreeRTOS_sys_clk sys_clk (
		.clk        (clock_sys_clk_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	FreeRTOS_timer_0 timer_0 (
		.clk        (clock_sys_clk_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	FreeRTOS_timer_0 timer_1 (
		.clk        (clock_sys_clk_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	FreeRTOS_timer_0 timer_2 (
		.clk        (clock_sys_clk_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_2_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_2_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_2_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_2_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_2_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver4_irq)                 //   irq.irq
	);

	FreeRTOS_mm_interconnect_0 mm_interconnect_0 (
		.clock_sys_clk_clk                              (clock_sys_clk_clk),                                           //                            clock_sys_clk.clk
		.FreeRTOSNios_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // FreeRTOSNios_reset_reset_bridge_in_reset.reset
		.FreeRTOSNios_data_master_address               (freertosnios_data_master_address),                            //                 FreeRTOSNios_data_master.address
		.FreeRTOSNios_data_master_waitrequest           (freertosnios_data_master_waitrequest),                        //                                         .waitrequest
		.FreeRTOSNios_data_master_byteenable            (freertosnios_data_master_byteenable),                         //                                         .byteenable
		.FreeRTOSNios_data_master_read                  (freertosnios_data_master_read),                               //                                         .read
		.FreeRTOSNios_data_master_readdata              (freertosnios_data_master_readdata),                           //                                         .readdata
		.FreeRTOSNios_data_master_readdatavalid         (freertosnios_data_master_readdatavalid),                      //                                         .readdatavalid
		.FreeRTOSNios_data_master_write                 (freertosnios_data_master_write),                              //                                         .write
		.FreeRTOSNios_data_master_writedata             (freertosnios_data_master_writedata),                          //                                         .writedata
		.FreeRTOSNios_data_master_debugaccess           (freertosnios_data_master_debugaccess),                        //                                         .debugaccess
		.FreeRTOSNios_instruction_master_address        (freertosnios_instruction_master_address),                     //          FreeRTOSNios_instruction_master.address
		.FreeRTOSNios_instruction_master_waitrequest    (freertosnios_instruction_master_waitrequest),                 //                                         .waitrequest
		.FreeRTOSNios_instruction_master_read           (freertosnios_instruction_master_read),                        //                                         .read
		.FreeRTOSNios_instruction_master_readdata       (freertosnios_instruction_master_readdata),                    //                                         .readdata
		.FreeRTOSNios_instruction_master_readdatavalid  (freertosnios_instruction_master_readdatavalid),               //                                         .readdatavalid
		.FreeRTOSNios_debug_mem_slave_address           (mm_interconnect_0_freertosnios_debug_mem_slave_address),      //             FreeRTOSNios_debug_mem_slave.address
		.FreeRTOSNios_debug_mem_slave_write             (mm_interconnect_0_freertosnios_debug_mem_slave_write),        //                                         .write
		.FreeRTOSNios_debug_mem_slave_read              (mm_interconnect_0_freertosnios_debug_mem_slave_read),         //                                         .read
		.FreeRTOSNios_debug_mem_slave_readdata          (mm_interconnect_0_freertosnios_debug_mem_slave_readdata),     //                                         .readdata
		.FreeRTOSNios_debug_mem_slave_writedata         (mm_interconnect_0_freertosnios_debug_mem_slave_writedata),    //                                         .writedata
		.FreeRTOSNios_debug_mem_slave_byteenable        (mm_interconnect_0_freertosnios_debug_mem_slave_byteenable),   //                                         .byteenable
		.FreeRTOSNios_debug_mem_slave_waitrequest       (mm_interconnect_0_freertosnios_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.FreeRTOSNios_debug_mem_slave_debugaccess       (mm_interconnect_0_freertosnios_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.Hex_0_avalon_slave_0_address                   (mm_interconnect_0_hex_0_avalon_slave_0_address),              //                     Hex_0_avalon_slave_0.address
		.Hex_0_avalon_slave_0_write                     (mm_interconnect_0_hex_0_avalon_slave_0_write),                //                                         .write
		.Hex_0_avalon_slave_0_readdata                  (mm_interconnect_0_hex_0_avalon_slave_0_readdata),             //                                         .readdata
		.Hex_0_avalon_slave_0_writedata                 (mm_interconnect_0_hex_0_avalon_slave_0_writedata),            //                                         .writedata
		.Hex_0_avalon_slave_0_chipselect                (mm_interconnect_0_hex_0_avalon_slave_0_chipselect),           //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.Piezo_0_avalon_slave_0_address                 (mm_interconnect_0_piezo_0_avalon_slave_0_address),            //                   Piezo_0_avalon_slave_0.address
		.Piezo_0_avalon_slave_0_write                   (mm_interconnect_0_piezo_0_avalon_slave_0_write),              //                                         .write
		.Piezo_0_avalon_slave_0_readdata                (mm_interconnect_0_piezo_0_avalon_slave_0_readdata),           //                                         .readdata
		.Piezo_0_avalon_slave_0_writedata               (mm_interconnect_0_piezo_0_avalon_slave_0_writedata),          //                                         .writedata
		.Piezo_0_avalon_slave_0_chipselect              (mm_interconnect_0_piezo_0_avalon_slave_0_chipselect),         //                                         .chipselect
		.sdram_s1_address                               (mm_interconnect_0_sdram_s1_address),                          //                                 sdram_s1.address
		.sdram_s1_write                                 (mm_interconnect_0_sdram_s1_write),                            //                                         .write
		.sdram_s1_read                                  (mm_interconnect_0_sdram_s1_read),                             //                                         .read
		.sdram_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                         //                                         .readdata
		.sdram_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                        //                                         .writedata
		.sdram_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                       //                                         .byteenable
		.sdram_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                         .readdatavalid
		.sdram_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),                      //                                         .waitrequest
		.sdram_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect),                       //                                         .chipselect
		.Servo_0_avalon_slave_0_address                 (mm_interconnect_0_servo_0_avalon_slave_0_address),            //                   Servo_0_avalon_slave_0.address
		.Servo_0_avalon_slave_0_write                   (mm_interconnect_0_servo_0_avalon_slave_0_write),              //                                         .write
		.Servo_0_avalon_slave_0_readdata                (mm_interconnect_0_servo_0_avalon_slave_0_readdata),           //                                         .readdata
		.Servo_0_avalon_slave_0_writedata               (mm_interconnect_0_servo_0_avalon_slave_0_writedata),          //                                         .writedata
		.Servo_0_avalon_slave_0_chipselect              (mm_interconnect_0_servo_0_avalon_slave_0_chipselect),         //                                         .chipselect
		.Servo_1_avalon_slave_0_address                 (mm_interconnect_0_servo_1_avalon_slave_0_address),            //                   Servo_1_avalon_slave_0.address
		.Servo_1_avalon_slave_0_write                   (mm_interconnect_0_servo_1_avalon_slave_0_write),              //                                         .write
		.Servo_1_avalon_slave_0_readdata                (mm_interconnect_0_servo_1_avalon_slave_0_readdata),           //                                         .readdata
		.Servo_1_avalon_slave_0_writedata               (mm_interconnect_0_servo_1_avalon_slave_0_writedata),          //                                         .writedata
		.Servo_1_avalon_slave_0_chipselect              (mm_interconnect_0_servo_1_avalon_slave_0_chipselect),         //                                         .chipselect
		.SW_0_avalon_slave_0_address                    (mm_interconnect_0_sw_0_avalon_slave_0_address),               //                      SW_0_avalon_slave_0.address
		.SW_0_avalon_slave_0_readdata                   (mm_interconnect_0_sw_0_avalon_slave_0_readdata),              //                                         .readdata
		.sys_clk_s1_address                             (mm_interconnect_0_sys_clk_s1_address),                        //                               sys_clk_s1.address
		.sys_clk_s1_write                               (mm_interconnect_0_sys_clk_s1_write),                          //                                         .write
		.sys_clk_s1_readdata                            (mm_interconnect_0_sys_clk_s1_readdata),                       //                                         .readdata
		.sys_clk_s1_writedata                           (mm_interconnect_0_sys_clk_s1_writedata),                      //                                         .writedata
		.sys_clk_s1_chipselect                          (mm_interconnect_0_sys_clk_s1_chipselect),                     //                                         .chipselect
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                        //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                          //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                       //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                      //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect),                     //                                         .chipselect
		.timer_1_s1_address                             (mm_interconnect_0_timer_1_s1_address),                        //                               timer_1_s1.address
		.timer_1_s1_write                               (mm_interconnect_0_timer_1_s1_write),                          //                                         .write
		.timer_1_s1_readdata                            (mm_interconnect_0_timer_1_s1_readdata),                       //                                         .readdata
		.timer_1_s1_writedata                           (mm_interconnect_0_timer_1_s1_writedata),                      //                                         .writedata
		.timer_1_s1_chipselect                          (mm_interconnect_0_timer_1_s1_chipselect),                     //                                         .chipselect
		.timer_2_s1_address                             (mm_interconnect_0_timer_2_s1_address),                        //                               timer_2_s1.address
		.timer_2_s1_write                               (mm_interconnect_0_timer_2_s1_write),                          //                                         .write
		.timer_2_s1_readdata                            (mm_interconnect_0_timer_2_s1_readdata),                       //                                         .readdata
		.timer_2_s1_writedata                           (mm_interconnect_0_timer_2_s1_writedata),                      //                                         .writedata
		.timer_2_s1_chipselect                          (mm_interconnect_0_timer_2_s1_chipselect)                      //                                         .chipselect
	);

	FreeRTOS_irq_mapper irq_mapper (
		.clk           (clock_sys_clk_clk),              //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (freertosnios_irq_irq)            //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (freertosnios_debug_reset_request_reset), // reset_in0.reset
		.clk            (clock_sys_clk_clk),                      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
