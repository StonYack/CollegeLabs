// Midterm.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module Midterm (
		input  wire        clk_clk,          //        clk.clk
		output wire [6:0]  hex_0_export,     //      hex_0.export
		output wire [6:0]  hex_1_export,     //      hex_1.export
		output wire [6:0]  hex_2_export,     //      hex_2.export
		output wire [6:0]  hex_3_export,     //      hex_3.export
		output wire [6:0]  hex_4_export,     //      hex_4.export
		output wire [6:0]  hex_5_export,     //      hex_5.export
		input  wire [3:0]  keys_export,      //       keys.export
		output wire [9:0]  leds_export,      //       leds.export
		output wire        sdram_clk_clk,    //  sdram_clk.clk
		output wire [12:0] sdram_wire_addr,  // sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,    //           .ba
		output wire        sdram_wire_cas_n, //           .cas_n
		output wire        sdram_wire_cke,   //           .cke
		output wire        sdram_wire_cs_n,  //           .cs_n
		inout  wire [15:0] sdram_wire_dq,    //           .dq
		output wire [1:0]  sdram_wire_dqm,   //           .dqm
		output wire        sdram_wire_ras_n, //           .ras_n
		output wire        sdram_wire_we_n,  //           .we_n
		input  wire [9:0]  sw_export         //         sw.export
	);

	wire         clock_sys_clk_clk;                                           // clock:sys_clk_clk -> [Hex_0:clk, Hex_1:clk, Hex_2:clk, Hex_3:clk, Hex_4:clk, Hex_5:clk, Keys:clk, Leds:clk, Midterm:clk, Switches:clk, irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:clock_sys_clk_clk, rst_controller:clk, sdram:clk, sys_clk:clk]
	wire         midterm_debug_reset_request_reset;                           // Midterm:debug_reset_request -> [clock:ref_reset_reset, rst_controller:reset_in0]
	wire  [31:0] midterm_data_master_readdata;                                // mm_interconnect_0:Midterm_data_master_readdata -> Midterm:d_readdata
	wire         midterm_data_master_waitrequest;                             // mm_interconnect_0:Midterm_data_master_waitrequest -> Midterm:d_waitrequest
	wire         midterm_data_master_debugaccess;                             // Midterm:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Midterm_data_master_debugaccess
	wire  [27:0] midterm_data_master_address;                                 // Midterm:d_address -> mm_interconnect_0:Midterm_data_master_address
	wire   [3:0] midterm_data_master_byteenable;                              // Midterm:d_byteenable -> mm_interconnect_0:Midterm_data_master_byteenable
	wire         midterm_data_master_read;                                    // Midterm:d_read -> mm_interconnect_0:Midterm_data_master_read
	wire         midterm_data_master_readdatavalid;                           // mm_interconnect_0:Midterm_data_master_readdatavalid -> Midterm:d_readdatavalid
	wire         midterm_data_master_write;                                   // Midterm:d_write -> mm_interconnect_0:Midterm_data_master_write
	wire  [31:0] midterm_data_master_writedata;                               // Midterm:d_writedata -> mm_interconnect_0:Midterm_data_master_writedata
	wire  [31:0] midterm_instruction_master_readdata;                         // mm_interconnect_0:Midterm_instruction_master_readdata -> Midterm:i_readdata
	wire         midterm_instruction_master_waitrequest;                      // mm_interconnect_0:Midterm_instruction_master_waitrequest -> Midterm:i_waitrequest
	wire  [26:0] midterm_instruction_master_address;                          // Midterm:i_address -> mm_interconnect_0:Midterm_instruction_master_address
	wire         midterm_instruction_master_read;                             // Midterm:i_read -> mm_interconnect_0:Midterm_instruction_master_read
	wire         midterm_instruction_master_readdatavalid;                    // mm_interconnect_0:Midterm_instruction_master_readdatavalid -> Midterm:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_switches_avalon_slave_0_readdata;          // Switches:readdata -> mm_interconnect_0:Switches_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_switches_avalon_slave_0_address;           // mm_interconnect_0:Switches_avalon_slave_0_address -> Switches:address
	wire         mm_interconnect_0_hex_0_avalon_slave_0_chipselect;           // mm_interconnect_0:Hex_0_avalon_slave_0_chipselect -> Hex_0:chipselect
	wire  [31:0] mm_interconnect_0_hex_0_avalon_slave_0_readdata;             // Hex_0:readdata -> mm_interconnect_0:Hex_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_hex_0_avalon_slave_0_address;              // mm_interconnect_0:Hex_0_avalon_slave_0_address -> Hex_0:address
	wire         mm_interconnect_0_hex_0_avalon_slave_0_write;                // mm_interconnect_0:Hex_0_avalon_slave_0_write -> Hex_0:write_n
	wire  [31:0] mm_interconnect_0_hex_0_avalon_slave_0_writedata;            // mm_interconnect_0:Hex_0_avalon_slave_0_writedata -> Hex_0:writedata
	wire         mm_interconnect_0_hex_1_avalon_slave_0_chipselect;           // mm_interconnect_0:Hex_1_avalon_slave_0_chipselect -> Hex_1:chipselect
	wire  [31:0] mm_interconnect_0_hex_1_avalon_slave_0_readdata;             // Hex_1:readdata -> mm_interconnect_0:Hex_1_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_hex_1_avalon_slave_0_address;              // mm_interconnect_0:Hex_1_avalon_slave_0_address -> Hex_1:address
	wire         mm_interconnect_0_hex_1_avalon_slave_0_write;                // mm_interconnect_0:Hex_1_avalon_slave_0_write -> Hex_1:write_n
	wire  [31:0] mm_interconnect_0_hex_1_avalon_slave_0_writedata;            // mm_interconnect_0:Hex_1_avalon_slave_0_writedata -> Hex_1:writedata
	wire         mm_interconnect_0_hex_2_avalon_slave_0_chipselect;           // mm_interconnect_0:Hex_2_avalon_slave_0_chipselect -> Hex_2:chipselect
	wire  [31:0] mm_interconnect_0_hex_2_avalon_slave_0_readdata;             // Hex_2:readdata -> mm_interconnect_0:Hex_2_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_hex_2_avalon_slave_0_address;              // mm_interconnect_0:Hex_2_avalon_slave_0_address -> Hex_2:address
	wire         mm_interconnect_0_hex_2_avalon_slave_0_write;                // mm_interconnect_0:Hex_2_avalon_slave_0_write -> Hex_2:write_n
	wire  [31:0] mm_interconnect_0_hex_2_avalon_slave_0_writedata;            // mm_interconnect_0:Hex_2_avalon_slave_0_writedata -> Hex_2:writedata
	wire         mm_interconnect_0_hex_3_avalon_slave_0_chipselect;           // mm_interconnect_0:Hex_3_avalon_slave_0_chipselect -> Hex_3:chipselect
	wire  [31:0] mm_interconnect_0_hex_3_avalon_slave_0_readdata;             // Hex_3:readdata -> mm_interconnect_0:Hex_3_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_hex_3_avalon_slave_0_address;              // mm_interconnect_0:Hex_3_avalon_slave_0_address -> Hex_3:address
	wire         mm_interconnect_0_hex_3_avalon_slave_0_write;                // mm_interconnect_0:Hex_3_avalon_slave_0_write -> Hex_3:write_n
	wire  [31:0] mm_interconnect_0_hex_3_avalon_slave_0_writedata;            // mm_interconnect_0:Hex_3_avalon_slave_0_writedata -> Hex_3:writedata
	wire         mm_interconnect_0_hex_4_avalon_slave_0_chipselect;           // mm_interconnect_0:Hex_4_avalon_slave_0_chipselect -> Hex_4:chipselect
	wire  [31:0] mm_interconnect_0_hex_4_avalon_slave_0_readdata;             // Hex_4:readdata -> mm_interconnect_0:Hex_4_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_hex_4_avalon_slave_0_address;              // mm_interconnect_0:Hex_4_avalon_slave_0_address -> Hex_4:address
	wire         mm_interconnect_0_hex_4_avalon_slave_0_write;                // mm_interconnect_0:Hex_4_avalon_slave_0_write -> Hex_4:write_n
	wire  [31:0] mm_interconnect_0_hex_4_avalon_slave_0_writedata;            // mm_interconnect_0:Hex_4_avalon_slave_0_writedata -> Hex_4:writedata
	wire         mm_interconnect_0_hex_5_avalon_slave_0_chipselect;           // mm_interconnect_0:Hex_5_avalon_slave_0_chipselect -> Hex_5:chipselect
	wire  [31:0] mm_interconnect_0_hex_5_avalon_slave_0_readdata;             // Hex_5:readdata -> mm_interconnect_0:Hex_5_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_hex_5_avalon_slave_0_address;              // mm_interconnect_0:Hex_5_avalon_slave_0_address -> Hex_5:address
	wire         mm_interconnect_0_hex_5_avalon_slave_0_write;                // mm_interconnect_0:Hex_5_avalon_slave_0_write -> Hex_5:write_n
	wire  [31:0] mm_interconnect_0_hex_5_avalon_slave_0_writedata;            // mm_interconnect_0:Hex_5_avalon_slave_0_writedata -> Hex_5:writedata
	wire  [31:0] mm_interconnect_0_keys_avalon_slave_0_readdata;              // Keys:readdata -> mm_interconnect_0:Keys_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_keys_avalon_slave_0_address;               // mm_interconnect_0:Keys_avalon_slave_0_address -> Keys:address
	wire         mm_interconnect_0_leds_avalon_slave_0_chipselect;            // mm_interconnect_0:Leds_avalon_slave_0_chipselect -> Leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_avalon_slave_0_readdata;              // Leds:readdata -> mm_interconnect_0:Leds_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_leds_avalon_slave_0_address;               // mm_interconnect_0:Leds_avalon_slave_0_address -> Leds:address
	wire         mm_interconnect_0_leds_avalon_slave_0_write;                 // mm_interconnect_0:Leds_avalon_slave_0_write -> Leds:write_n
	wire  [31:0] mm_interconnect_0_leds_avalon_slave_0_writedata;             // mm_interconnect_0:Leds_avalon_slave_0_writedata -> Leds:writedata
	wire  [31:0] mm_interconnect_0_midterm_debug_mem_slave_readdata;          // Midterm:debug_mem_slave_readdata -> mm_interconnect_0:Midterm_debug_mem_slave_readdata
	wire         mm_interconnect_0_midterm_debug_mem_slave_waitrequest;       // Midterm:debug_mem_slave_waitrequest -> mm_interconnect_0:Midterm_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_midterm_debug_mem_slave_debugaccess;       // mm_interconnect_0:Midterm_debug_mem_slave_debugaccess -> Midterm:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_midterm_debug_mem_slave_address;           // mm_interconnect_0:Midterm_debug_mem_slave_address -> Midterm:debug_mem_slave_address
	wire         mm_interconnect_0_midterm_debug_mem_slave_read;              // mm_interconnect_0:Midterm_debug_mem_slave_read -> Midterm:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_midterm_debug_mem_slave_byteenable;        // mm_interconnect_0:Midterm_debug_mem_slave_byteenable -> Midterm:debug_mem_slave_byteenable
	wire         mm_interconnect_0_midterm_debug_mem_slave_write;             // mm_interconnect_0:Midterm_debug_mem_slave_write -> Midterm:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_midterm_debug_mem_slave_writedata;         // mm_interconnect_0:Midterm_debug_mem_slave_writedata -> Midterm:debug_mem_slave_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                         // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_sys_clk_s1_chipselect;                     // mm_interconnect_0:sys_clk_s1_chipselect -> sys_clk:chipselect
	wire  [15:0] mm_interconnect_0_sys_clk_s1_readdata;                       // sys_clk:readdata -> mm_interconnect_0:sys_clk_s1_readdata
	wire   [2:0] mm_interconnect_0_sys_clk_s1_address;                        // mm_interconnect_0:sys_clk_s1_address -> sys_clk:address
	wire         mm_interconnect_0_sys_clk_s1_write;                          // mm_interconnect_0:sys_clk_s1_write -> sys_clk:write_n
	wire  [15:0] mm_interconnect_0_sys_clk_s1_writedata;                      // mm_interconnect_0:sys_clk_s1_writedata -> sys_clk:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // sys_clk:irq -> irq_mapper:receiver1_irq
	wire  [31:0] midterm_irq_irq;                                             // irq_mapper:sender_irq -> Midterm:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [Hex_0:reset_n, Hex_1:reset_n, Hex_2:reset_n, Hex_3:reset_n, Hex_4:reset_n, Hex_5:reset_n, Keys:reset_n, Leds:reset_n, Midterm:reset_n, Switches:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:Midterm_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sdram:reset_n, sys_clk:reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [Midterm:reset_req, rst_translator:reset_req_in]

	My_Hex hex_0 (
		.address    (mm_interconnect_0_hex_0_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_hex_0_avalon_slave_0_chipselect), //               .chipselect
		.write_n    (~mm_interconnect_0_hex_0_avalon_slave_0_write),     //               .write_n
		.writedata  (mm_interconnect_0_hex_0_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_hex_0_avalon_slave_0_readdata),   //               .readdata
		.clk        (clock_sys_clk_clk),                                 //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //          reset.reset_n
		.out_port   (hex_0_export)                                       //    conduit_end.export
	);

	My_Hex hex_1 (
		.address    (mm_interconnect_0_hex_1_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_hex_1_avalon_slave_0_chipselect), //               .chipselect
		.write_n    (~mm_interconnect_0_hex_1_avalon_slave_0_write),     //               .write_n
		.writedata  (mm_interconnect_0_hex_1_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_hex_1_avalon_slave_0_readdata),   //               .readdata
		.clk        (clock_sys_clk_clk),                                 //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //          reset.reset_n
		.out_port   (hex_1_export)                                       //    conduit_end.export
	);

	My_Hex hex_2 (
		.address    (mm_interconnect_0_hex_2_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_hex_2_avalon_slave_0_chipselect), //               .chipselect
		.write_n    (~mm_interconnect_0_hex_2_avalon_slave_0_write),     //               .write_n
		.writedata  (mm_interconnect_0_hex_2_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_hex_2_avalon_slave_0_readdata),   //               .readdata
		.clk        (clock_sys_clk_clk),                                 //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //          reset.reset_n
		.out_port   (hex_2_export)                                       //    conduit_end.export
	);

	My_Hex hex_3 (
		.address    (mm_interconnect_0_hex_3_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_hex_3_avalon_slave_0_chipselect), //               .chipselect
		.write_n    (~mm_interconnect_0_hex_3_avalon_slave_0_write),     //               .write_n
		.writedata  (mm_interconnect_0_hex_3_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_hex_3_avalon_slave_0_readdata),   //               .readdata
		.clk        (clock_sys_clk_clk),                                 //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //          reset.reset_n
		.out_port   (hex_3_export)                                       //    conduit_end.export
	);

	My_Hex hex_4 (
		.address    (mm_interconnect_0_hex_4_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_hex_4_avalon_slave_0_chipselect), //               .chipselect
		.write_n    (~mm_interconnect_0_hex_4_avalon_slave_0_write),     //               .write_n
		.writedata  (mm_interconnect_0_hex_4_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_hex_4_avalon_slave_0_readdata),   //               .readdata
		.clk        (clock_sys_clk_clk),                                 //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //          reset.reset_n
		.out_port   (hex_4_export)                                       //    conduit_end.export
	);

	My_Hex hex_5 (
		.address    (mm_interconnect_0_hex_5_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_hex_5_avalon_slave_0_chipselect), //               .chipselect
		.write_n    (~mm_interconnect_0_hex_5_avalon_slave_0_write),     //               .write_n
		.writedata  (mm_interconnect_0_hex_5_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_hex_5_avalon_slave_0_readdata),   //               .readdata
		.clk        (clock_sys_clk_clk),                                 //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //          reset.reset_n
		.out_port   (hex_5_export)                                       //    conduit_end.export
	);

	My_Key keys (
		.address  (mm_interconnect_0_keys_avalon_slave_0_address),  // avalon_slave_0.address
		.readdata (mm_interconnect_0_keys_avalon_slave_0_readdata), //               .readdata
		.clk      (clock_sys_clk_clk),                              //          clock.clk
		.reset_n  (~rst_controller_reset_out_reset),                //          reset.reset_n
		.Key_in   (keys_export)                                     //    conduit_end.export
	);

	My_Led leds (
		.address    (mm_interconnect_0_leds_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect (mm_interconnect_0_leds_avalon_slave_0_chipselect), //               .chipselect
		.write_n    (~mm_interconnect_0_leds_avalon_slave_0_write),     //               .write_n
		.writedata  (mm_interconnect_0_leds_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_leds_avalon_slave_0_readdata),   //               .readdata
		.clk        (clock_sys_clk_clk),                                //          clock.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //          reset.reset_n
		.out_port   (leds_export)                                       //    conduit_end.export
	);

	Midterm_Midterm midterm (
		.clk                                 (clock_sys_clk_clk),                                     //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                       //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                           (midterm_data_master_address),                           //               data_master.address
		.d_byteenable                        (midterm_data_master_byteenable),                        //                          .byteenable
		.d_read                              (midterm_data_master_read),                              //                          .read
		.d_readdata                          (midterm_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (midterm_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (midterm_data_master_write),                             //                          .write
		.d_writedata                         (midterm_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (midterm_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (midterm_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (midterm_instruction_master_address),                    //        instruction_master.address
		.i_read                              (midterm_instruction_master_read),                       //                          .read
		.i_readdata                          (midterm_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (midterm_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (midterm_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (midterm_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (midterm_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_midterm_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_midterm_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_midterm_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_midterm_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_midterm_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_midterm_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_midterm_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_midterm_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                       // custom_instruction_master.readra
	);

	My_SW switches (
		.address  (mm_interconnect_0_switches_avalon_slave_0_address),  // avalon_slave_0.address
		.readdata (mm_interconnect_0_switches_avalon_slave_0_readdata), //               .readdata
		.clk      (clock_sys_clk_clk),                                  //          clock.clk
		.reset_n  (~rst_controller_reset_out_reset),                    //          reset.reset_n
		.SW_in    (sw_export)                                           //    conduit_end.export
	);

	Midterm_clock clock (
		.ref_clk_clk        (clk_clk),                           //      ref_clk.clk
		.ref_reset_reset    (midterm_debug_reset_request_reset), //    ref_reset.reset
		.sys_clk_clk        (clock_sys_clk_clk),                 //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                     //    sdram_clk.clk
		.reset_source_reset ()                                   // reset_source.reset
	);

	Midterm_jtag_uart_0 jtag_uart_0 (
		.clk            (clock_sys_clk_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	Midterm_sdram sdram (
		.clk            (clock_sys_clk_clk),                        //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	Midterm_sys_clk sys_clk (
		.clk        (clock_sys_clk_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_sys_clk_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_clk_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_clk_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_clk_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_clk_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	Midterm_mm_interconnect_0 mm_interconnect_0 (
		.clock_sys_clk_clk                         (clock_sys_clk_clk),                                           //                       clock_sys_clk.clk
		.Midterm_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // Midterm_reset_reset_bridge_in_reset.reset
		.Midterm_data_master_address               (midterm_data_master_address),                                 //                 Midterm_data_master.address
		.Midterm_data_master_waitrequest           (midterm_data_master_waitrequest),                             //                                    .waitrequest
		.Midterm_data_master_byteenable            (midterm_data_master_byteenable),                              //                                    .byteenable
		.Midterm_data_master_read                  (midterm_data_master_read),                                    //                                    .read
		.Midterm_data_master_readdata              (midterm_data_master_readdata),                                //                                    .readdata
		.Midterm_data_master_readdatavalid         (midterm_data_master_readdatavalid),                           //                                    .readdatavalid
		.Midterm_data_master_write                 (midterm_data_master_write),                                   //                                    .write
		.Midterm_data_master_writedata             (midterm_data_master_writedata),                               //                                    .writedata
		.Midterm_data_master_debugaccess           (midterm_data_master_debugaccess),                             //                                    .debugaccess
		.Midterm_instruction_master_address        (midterm_instruction_master_address),                          //          Midterm_instruction_master.address
		.Midterm_instruction_master_waitrequest    (midterm_instruction_master_waitrequest),                      //                                    .waitrequest
		.Midterm_instruction_master_read           (midterm_instruction_master_read),                             //                                    .read
		.Midterm_instruction_master_readdata       (midterm_instruction_master_readdata),                         //                                    .readdata
		.Midterm_instruction_master_readdatavalid  (midterm_instruction_master_readdatavalid),                    //                                    .readdatavalid
		.Hex_0_avalon_slave_0_address              (mm_interconnect_0_hex_0_avalon_slave_0_address),              //                Hex_0_avalon_slave_0.address
		.Hex_0_avalon_slave_0_write                (mm_interconnect_0_hex_0_avalon_slave_0_write),                //                                    .write
		.Hex_0_avalon_slave_0_readdata             (mm_interconnect_0_hex_0_avalon_slave_0_readdata),             //                                    .readdata
		.Hex_0_avalon_slave_0_writedata            (mm_interconnect_0_hex_0_avalon_slave_0_writedata),            //                                    .writedata
		.Hex_0_avalon_slave_0_chipselect           (mm_interconnect_0_hex_0_avalon_slave_0_chipselect),           //                                    .chipselect
		.Hex_1_avalon_slave_0_address              (mm_interconnect_0_hex_1_avalon_slave_0_address),              //                Hex_1_avalon_slave_0.address
		.Hex_1_avalon_slave_0_write                (mm_interconnect_0_hex_1_avalon_slave_0_write),                //                                    .write
		.Hex_1_avalon_slave_0_readdata             (mm_interconnect_0_hex_1_avalon_slave_0_readdata),             //                                    .readdata
		.Hex_1_avalon_slave_0_writedata            (mm_interconnect_0_hex_1_avalon_slave_0_writedata),            //                                    .writedata
		.Hex_1_avalon_slave_0_chipselect           (mm_interconnect_0_hex_1_avalon_slave_0_chipselect),           //                                    .chipselect
		.Hex_2_avalon_slave_0_address              (mm_interconnect_0_hex_2_avalon_slave_0_address),              //                Hex_2_avalon_slave_0.address
		.Hex_2_avalon_slave_0_write                (mm_interconnect_0_hex_2_avalon_slave_0_write),                //                                    .write
		.Hex_2_avalon_slave_0_readdata             (mm_interconnect_0_hex_2_avalon_slave_0_readdata),             //                                    .readdata
		.Hex_2_avalon_slave_0_writedata            (mm_interconnect_0_hex_2_avalon_slave_0_writedata),            //                                    .writedata
		.Hex_2_avalon_slave_0_chipselect           (mm_interconnect_0_hex_2_avalon_slave_0_chipselect),           //                                    .chipselect
		.Hex_3_avalon_slave_0_address              (mm_interconnect_0_hex_3_avalon_slave_0_address),              //                Hex_3_avalon_slave_0.address
		.Hex_3_avalon_slave_0_write                (mm_interconnect_0_hex_3_avalon_slave_0_write),                //                                    .write
		.Hex_3_avalon_slave_0_readdata             (mm_interconnect_0_hex_3_avalon_slave_0_readdata),             //                                    .readdata
		.Hex_3_avalon_slave_0_writedata            (mm_interconnect_0_hex_3_avalon_slave_0_writedata),            //                                    .writedata
		.Hex_3_avalon_slave_0_chipselect           (mm_interconnect_0_hex_3_avalon_slave_0_chipselect),           //                                    .chipselect
		.Hex_4_avalon_slave_0_address              (mm_interconnect_0_hex_4_avalon_slave_0_address),              //                Hex_4_avalon_slave_0.address
		.Hex_4_avalon_slave_0_write                (mm_interconnect_0_hex_4_avalon_slave_0_write),                //                                    .write
		.Hex_4_avalon_slave_0_readdata             (mm_interconnect_0_hex_4_avalon_slave_0_readdata),             //                                    .readdata
		.Hex_4_avalon_slave_0_writedata            (mm_interconnect_0_hex_4_avalon_slave_0_writedata),            //                                    .writedata
		.Hex_4_avalon_slave_0_chipselect           (mm_interconnect_0_hex_4_avalon_slave_0_chipselect),           //                                    .chipselect
		.Hex_5_avalon_slave_0_address              (mm_interconnect_0_hex_5_avalon_slave_0_address),              //                Hex_5_avalon_slave_0.address
		.Hex_5_avalon_slave_0_write                (mm_interconnect_0_hex_5_avalon_slave_0_write),                //                                    .write
		.Hex_5_avalon_slave_0_readdata             (mm_interconnect_0_hex_5_avalon_slave_0_readdata),             //                                    .readdata
		.Hex_5_avalon_slave_0_writedata            (mm_interconnect_0_hex_5_avalon_slave_0_writedata),            //                                    .writedata
		.Hex_5_avalon_slave_0_chipselect           (mm_interconnect_0_hex_5_avalon_slave_0_chipselect),           //                                    .chipselect
		.jtag_uart_0_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //       jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                    .write
		.jtag_uart_0_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                    .read
		.jtag_uart_0_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                    .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                    .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                    .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                    .chipselect
		.Keys_avalon_slave_0_address               (mm_interconnect_0_keys_avalon_slave_0_address),               //                 Keys_avalon_slave_0.address
		.Keys_avalon_slave_0_readdata              (mm_interconnect_0_keys_avalon_slave_0_readdata),              //                                    .readdata
		.Leds_avalon_slave_0_address               (mm_interconnect_0_leds_avalon_slave_0_address),               //                 Leds_avalon_slave_0.address
		.Leds_avalon_slave_0_write                 (mm_interconnect_0_leds_avalon_slave_0_write),                 //                                    .write
		.Leds_avalon_slave_0_readdata              (mm_interconnect_0_leds_avalon_slave_0_readdata),              //                                    .readdata
		.Leds_avalon_slave_0_writedata             (mm_interconnect_0_leds_avalon_slave_0_writedata),             //                                    .writedata
		.Leds_avalon_slave_0_chipselect            (mm_interconnect_0_leds_avalon_slave_0_chipselect),            //                                    .chipselect
		.Midterm_debug_mem_slave_address           (mm_interconnect_0_midterm_debug_mem_slave_address),           //             Midterm_debug_mem_slave.address
		.Midterm_debug_mem_slave_write             (mm_interconnect_0_midterm_debug_mem_slave_write),             //                                    .write
		.Midterm_debug_mem_slave_read              (mm_interconnect_0_midterm_debug_mem_slave_read),              //                                    .read
		.Midterm_debug_mem_slave_readdata          (mm_interconnect_0_midterm_debug_mem_slave_readdata),          //                                    .readdata
		.Midterm_debug_mem_slave_writedata         (mm_interconnect_0_midterm_debug_mem_slave_writedata),         //                                    .writedata
		.Midterm_debug_mem_slave_byteenable        (mm_interconnect_0_midterm_debug_mem_slave_byteenable),        //                                    .byteenable
		.Midterm_debug_mem_slave_waitrequest       (mm_interconnect_0_midterm_debug_mem_slave_waitrequest),       //                                    .waitrequest
		.Midterm_debug_mem_slave_debugaccess       (mm_interconnect_0_midterm_debug_mem_slave_debugaccess),       //                                    .debugaccess
		.sdram_s1_address                          (mm_interconnect_0_sdram_s1_address),                          //                            sdram_s1.address
		.sdram_s1_write                            (mm_interconnect_0_sdram_s1_write),                            //                                    .write
		.sdram_s1_read                             (mm_interconnect_0_sdram_s1_read),                             //                                    .read
		.sdram_s1_readdata                         (mm_interconnect_0_sdram_s1_readdata),                         //                                    .readdata
		.sdram_s1_writedata                        (mm_interconnect_0_sdram_s1_writedata),                        //                                    .writedata
		.sdram_s1_byteenable                       (mm_interconnect_0_sdram_s1_byteenable),                       //                                    .byteenable
		.sdram_s1_readdatavalid                    (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                    .readdatavalid
		.sdram_s1_waitrequest                      (mm_interconnect_0_sdram_s1_waitrequest),                      //                                    .waitrequest
		.sdram_s1_chipselect                       (mm_interconnect_0_sdram_s1_chipselect),                       //                                    .chipselect
		.Switches_avalon_slave_0_address           (mm_interconnect_0_switches_avalon_slave_0_address),           //             Switches_avalon_slave_0.address
		.Switches_avalon_slave_0_readdata          (mm_interconnect_0_switches_avalon_slave_0_readdata),          //                                    .readdata
		.sys_clk_s1_address                        (mm_interconnect_0_sys_clk_s1_address),                        //                          sys_clk_s1.address
		.sys_clk_s1_write                          (mm_interconnect_0_sys_clk_s1_write),                          //                                    .write
		.sys_clk_s1_readdata                       (mm_interconnect_0_sys_clk_s1_readdata),                       //                                    .readdata
		.sys_clk_s1_writedata                      (mm_interconnect_0_sys_clk_s1_writedata),                      //                                    .writedata
		.sys_clk_s1_chipselect                     (mm_interconnect_0_sys_clk_s1_chipselect)                      //                                    .chipselect
	);

	Midterm_irq_mapper irq_mapper (
		.clk           (clock_sys_clk_clk),              //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (midterm_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (midterm_debug_reset_request_reset),  // reset_in0.reset
		.clk            (clock_sys_clk_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
