
module Lab3Nios (
	clk_clk,
	hex_export,
	switches_export);	

	input		clk_clk;
	output	[20:0]	hex_export;
	input	[9:0]	switches_export;
endmodule
